LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY busMux_encoder IS
PORT(
	r00_out, r01_out, r02_out, r03_out,
	r04_out, r05_out, r06_out, r07_out,
	r08_out, r09_out, r10_out, r11_out,
	r12_out, r13_out, r14_out, r15_out,
	hi_out, lo_out, z_hi_out, z_lo_out,
	PC_out, MDR_out, port_out, c_out	: IN std_logic;
	s_out	:	OUT std_logic_vector(4 downto 0)
);
END busMux_encoder;

ARCHITECTURE behavioural OF busMux_encoder IS
BEGIN
	s_out <= 	"00000" when (r00_out='1')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='0') else
					"00001" when (r00_out='0')and(r01_out='1')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='0') else
					"00010" when (r00_out='0')and(r01_out='0')and(r02_out='1')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='0') else
					"00011" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='1')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='0') else
					"00100" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='1')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='0') else
					"00101" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='1')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='0') else
					"00110" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='1')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='0') else
					"00111" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='1')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='0') else
					"01000" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='1')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='0') else
					"01001" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='1')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='0') else
					"01010" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='1')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='0') else
					"01011" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='1')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='0') else
					"01100" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='1')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='0') else
					"01101" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='1')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='0') else
					"01110" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='1')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='0') else
					"01111" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='1')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='0') else
					"10000" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='1')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='0') else
					"10001" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='1')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='0') else
					"10010" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='1')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='0') else
					"10011" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='1')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='0') else
					"10100" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='1')and(MDR_out='0')and(port_out='0')and(c_out='0') else
					"10101" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='1')and(port_out='0')and(c_out='0') else
					"10110" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='1')and(c_out='0') else
					"10111" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='1') else
					"11110" when (r00_out='0')and(r01_out='0')and(r02_out='0')and(r03_out='0')and(r04_out='0')and(r05_out='0')and(r06_out='0')and(r07_out='0')and(r08_out='0')and(r09_out='0')and(r10_out='0')and(r11_out='0')and(r12_out='0')and(r13_out='0')and(r14_out='0')and(r15_out='0')and(hi_out='0')and(lo_out='0')and(z_hi_out='0')and(z_lo_out='0')and(PC_out='0')and(MDR_out='0')and(port_out='0')and(c_out='1') else
					--^ signal for no input
					"11111";
END behavioural;