LIBRARY IEEE;
USE ieee.std_logic_1164.all;

ENTITY cpu_codyale_ph3_tb IS
END ENTITY;

ARCHITECTURE behavioural OF cpu_codyale_ph3_tb IS 
COMPONENT cpu_codyale
	PORT(
	);
END COMPONENT;

BEGIN
	clk_process :PROCESS
	BEGIN
	END PROCESS;
	
	tb : PROCESS
	BEGIN
	END PROCESS;
END;